`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/09/04 13:37:57
// Design Name: 
// Module Name: CPU_test
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module CPU_test_tb();
    reg clk, rst, go;
//    wire [7:0] SEG;   // 7��������������͵�ƽ��Ч
//    wire [7:0] AN;    // 7�������Ƭѡ�źţ��͵�ƽ��Ч;
//    wire IRAin,IRBin,IRCin;
//    wire [15:0] circles;
//    wire [1:0] IntNo,clrNo;
//    wire uret,INT,IE;
//    wire [31:0] IntAddr;
//    wire [31:0] LedData, IR, ALU_result_F,AinF, BinF, FR1out,FR2out,FRDin,PCout;
//    wire Jal,Jalr,BJMP,clk_n,halt,ecall;
//    wire [4:0] ALU_OP_2,FR1in, FR2in,rd;
//    wire FMemtoReg,FMemWrite,ALU_Src,FRegWrite,itof,ftoi,RegWrite,auipc;
//    wire [31:0] Result,Memin_sb_ext,Memout,R2out,ALU_result1;
//    wire [7:0] Memin_sb;
    reg [25087:0] InputData;
    wire done;
    wire [31:0] Res;
      
    initial begin
        clk=0;
        rst=1;
        go=0;
        InputData[31:0] = 32'h00000000;
        InputData[63:32] = 32'h00000000;
        InputData[95:64] = 32'h00000000;
        InputData[127:96] = 32'h00000000;
        InputData[159:128] = 32'h00000000;
        InputData[191:160] = 32'h00000000;
        InputData[223:192] = 32'h00000000;
        InputData[255:224] = 32'h00000000;
        InputData[287:256] = 32'h00000000;
        InputData[319:288] = 32'h00000000;
        InputData[351:320] = 32'h00000000;
        InputData[383:352] = 32'h00000000;
        InputData[415:384] = 32'h00000000;
        InputData[447:416] = 32'h00000000;
        InputData[479:448] = 32'h00000000;
        InputData[511:480] = 32'h00000000;
        InputData[543:512] = 32'h00000000;
        InputData[575:544] = 32'h00000000;
        InputData[607:576] = 32'h00000000;
        InputData[639:608] = 32'h00000000;
        InputData[671:640] = 32'h00000000;
        InputData[703:672] = 32'h00000000;
        InputData[735:704] = 32'h00000000;
        InputData[767:736] = 32'h00000000;
        InputData[799:768] = 32'h00000000;
        InputData[831:800] = 32'h00000000;
        InputData[863:832] = 32'h00000000;
        InputData[895:864] = 32'h00000000;
        InputData[927:896] = 32'h00000000;
        InputData[959:928] = 32'h00000000;
        InputData[991:960] = 32'h00000000;
        InputData[1023:992] = 32'h00000000;
        InputData[1055:1024] = 32'h00000000;
        InputData[1087:1056] = 32'h00000000;
        InputData[1119:1088] = 32'h00000000;
        InputData[1151:1120] = 32'h00000000;
        InputData[1183:1152] = 32'h00000000;
        InputData[1215:1184] = 32'h00000000;
        InputData[1247:1216] = 32'h00000000;
        InputData[1279:1248] = 32'h00000000;
        InputData[1311:1280] = 32'h00000000;
        InputData[1343:1312] = 32'h00000000;
        InputData[1375:1344] = 32'h00000000;
        InputData[1407:1376] = 32'h00000000;
        InputData[1439:1408] = 32'h00000000;
        InputData[1471:1440] = 32'h00000000;
        InputData[1503:1472] = 32'h00000000;
        InputData[1535:1504] = 32'h00000000;
        InputData[1567:1536] = 32'h00000000;
        InputData[1599:1568] = 32'h00000000;
        InputData[1631:1600] = 32'h00000000;
        InputData[1663:1632] = 32'h00000000;
        InputData[1695:1664] = 32'h00000000;
        InputData[1727:1696] = 32'h00000000;
        InputData[1759:1728] = 32'h00000000;
        InputData[1791:1760] = 32'h00000000;
        InputData[1823:1792] = 32'h00000000;
        InputData[1855:1824] = 32'h00000000;
        InputData[1887:1856] = 32'h00000000;
        InputData[1919:1888] = 32'h00000000;
        InputData[1951:1920] = 32'h00000000;
        InputData[1983:1952] = 32'h00000000;
        InputData[2015:1984] = 32'h00000000;
        InputData[2047:2016] = 32'h00000000;
        InputData[2079:2048] = 32'h00000000;
        InputData[2111:2080] = 32'h00000000;
        InputData[2143:2112] = 32'h00000000;
        InputData[2175:2144] = 32'h00000000;
        InputData[2207:2176] = 32'h00000000;
        InputData[2239:2208] = 32'h00000000;
        InputData[2271:2240] = 32'h00000000;
        InputData[2303:2272] = 32'h00000000;
        InputData[2335:2304] = 32'h00000000;
        InputData[2367:2336] = 32'h00000000;
        InputData[2399:2368] = 32'h00000000;
        InputData[2431:2400] = 32'h00000000;
        InputData[2463:2432] = 32'h00000000;
        InputData[2495:2464] = 32'h00000000;
        InputData[2527:2496] = 32'h00000000;
        InputData[2559:2528] = 32'h00000000;
        InputData[2591:2560] = 32'h00000000;
        InputData[2623:2592] = 32'h00000000;
        InputData[2655:2624] = 32'h00000000;
        InputData[2687:2656] = 32'h00000000;
        InputData[2719:2688] = 32'h00000000;
        InputData[2751:2720] = 32'h00000000;
        InputData[2783:2752] = 32'h00000000;
        InputData[2815:2784] = 32'h00000000;
        InputData[2847:2816] = 32'h00000000;
        InputData[2879:2848] = 32'h00000000;
        InputData[2911:2880] = 32'h00000000;
        InputData[2943:2912] = 32'h00000000;
        InputData[2975:2944] = 32'h00000000;
        InputData[3007:2976] = 32'h00000000;
        InputData[3039:3008] = 32'h00000000;
        InputData[3071:3040] = 32'h00000000;
        InputData[3103:3072] = 32'h00000000;
        InputData[3135:3104] = 32'h00000000;
        InputData[3167:3136] = 32'h00000000;
        InputData[3199:3168] = 32'h00000000;
        InputData[3231:3200] = 32'h00000000;
        InputData[3263:3232] = 32'h00000000;
        InputData[3295:3264] = 32'h00000000;
        InputData[3327:3296] = 32'h00000000;
        InputData[3359:3328] = 32'h00000000;
        InputData[3391:3360] = 32'h00000000;
        InputData[3423:3392] = 32'h00000000;
        InputData[3455:3424] = 32'h00000000;
        InputData[3487:3456] = 32'h00000000;
        InputData[3519:3488] = 32'h00000000;
        InputData[3551:3520] = 32'h00000000;
        InputData[3583:3552] = 32'h00000000;
        InputData[3615:3584] = 32'h00000000;
        InputData[3647:3616] = 32'h00000000;
        InputData[3679:3648] = 32'h00000000;
        InputData[3711:3680] = 32'h00000000;
        InputData[3743:3712] = 32'h00000000;
        InputData[3775:3744] = 32'h00000000;
        InputData[3807:3776] = 32'h00000000;
        InputData[3839:3808] = 32'h00000000;
        InputData[3871:3840] = 32'h00000000;
        InputData[3903:3872] = 32'h00000000;
        InputData[3935:3904] = 32'h00000000;
        InputData[3967:3936] = 32'h3f800000;
        InputData[3999:3968] = 32'h3f800000;
        InputData[4031:4000] = 32'h3f800000;
        InputData[4063:4032] = 32'h00000000;
        InputData[4095:4064] = 32'h00000000;
        InputData[4127:4096] = 32'h00000000;
        InputData[4159:4128] = 32'h00000000;
        InputData[4191:4160] = 32'h00000000;
        InputData[4223:4192] = 32'h00000000;
        InputData[4255:4224] = 32'h00000000;
        InputData[4287:4256] = 32'h00000000;
        InputData[4319:4288] = 32'h00000000;
        InputData[4351:4320] = 32'h00000000;
        InputData[4383:4352] = 32'h00000000;
        InputData[4415:4384] = 32'h00000000;
        InputData[4447:4416] = 32'h00000000;
        InputData[4479:4448] = 32'h00000000;
        InputData[4511:4480] = 32'h00000000;
        InputData[4543:4512] = 32'h00000000;
        InputData[4575:4544] = 32'h00000000;
        InputData[4607:4576] = 32'h00000000;
        InputData[4639:4608] = 32'h00000000;
        InputData[4671:4640] = 32'h00000000;
        InputData[4703:4672] = 32'h00000000;
        InputData[4735:4704] = 32'h00000000;
        InputData[4767:4736] = 32'h00000000;
        InputData[4799:4768] = 32'h00000000;
        InputData[4831:4800] = 32'h00000000;
        InputData[4863:4832] = 32'h3f800000;
        InputData[4895:4864] = 32'h3f800000;
        InputData[4927:4896] = 32'h3f800000;
        InputData[4959:4928] = 32'h00000000;
        InputData[4991:4960] = 32'h00000000;
        InputData[5023:4992] = 32'h00000000;
        InputData[5055:5024] = 32'h00000000;
        InputData[5087:5056] = 32'h00000000;
        InputData[5119:5088] = 32'h00000000;
        InputData[5151:5120] = 32'h00000000;
        InputData[5183:5152] = 32'h3f800000;
        InputData[5215:5184] = 32'h3f800000;
        InputData[5247:5216] = 32'h00000000;
        InputData[5279:5248] = 32'h00000000;
        InputData[5311:5280] = 32'h00000000;
        InputData[5343:5312] = 32'h00000000;
        InputData[5375:5344] = 32'h00000000;
        InputData[5407:5376] = 32'h00000000;
        InputData[5439:5408] = 32'h00000000;
        InputData[5471:5440] = 32'h00000000;
        InputData[5503:5472] = 32'h00000000;
        InputData[5535:5504] = 32'h00000000;
        InputData[5567:5536] = 32'h00000000;
        InputData[5599:5568] = 32'h00000000;
        InputData[5631:5600] = 32'h00000000;
        InputData[5663:5632] = 32'h00000000;
        InputData[5695:5664] = 32'h00000000;
        InputData[5727:5696] = 32'h00000000;
        InputData[5759:5728] = 32'h3f800000;
        InputData[5791:5760] = 32'h3f800000;
        InputData[5823:5792] = 32'h3f800000;
        InputData[5855:5824] = 32'h00000000;
        InputData[5887:5856] = 32'h00000000;
        InputData[5919:5888] = 32'h00000000;
        InputData[5951:5920] = 32'h00000000;
        InputData[5983:5952] = 32'h00000000;
        InputData[6015:5984] = 32'h00000000;
        InputData[6047:6016] = 32'h3f800000;
        InputData[6079:6048] = 32'h3f800000;
        InputData[6111:6080] = 32'h3f800000;
        InputData[6143:6112] = 32'h00000000;
        InputData[6175:6144] = 32'h00000000;
        InputData[6207:6176] = 32'h00000000;
        InputData[6239:6208] = 32'h00000000;
        InputData[6271:6240] = 32'h00000000;
        InputData[6303:6272] = 32'h00000000;
        InputData[6335:6304] = 32'h00000000;
        InputData[6367:6336] = 32'h00000000;
        InputData[6399:6368] = 32'h00000000;
        InputData[6431:6400] = 32'h00000000;
        InputData[6463:6432] = 32'h00000000;
        InputData[6495:6464] = 32'h00000000;
        InputData[6527:6496] = 32'h00000000;
        InputData[6559:6528] = 32'h00000000;
        InputData[6591:6560] = 32'h00000000;
        InputData[6623:6592] = 32'h00000000;
        InputData[6655:6624] = 32'h3f800000;
        InputData[6687:6656] = 32'h3f800000;
        InputData[6719:6688] = 32'h3f800000;
        InputData[6751:6720] = 32'h00000000;
        InputData[6783:6752] = 32'h00000000;
        InputData[6815:6784] = 32'h00000000;
        InputData[6847:6816] = 32'h00000000;
        InputData[6879:6848] = 32'h00000000;
        InputData[6911:6880] = 32'h00000000;
        InputData[6943:6912] = 32'h3f800000;
        InputData[6975:6944] = 32'h3f800000;
        InputData[7007:6976] = 32'h3f800000;
        InputData[7039:7008] = 32'h00000000;
        InputData[7071:7040] = 32'h00000000;
        InputData[7103:7072] = 32'h00000000;
        InputData[7135:7104] = 32'h00000000;
        InputData[7167:7136] = 32'h00000000;
        InputData[7199:7168] = 32'h00000000;
        InputData[7231:7200] = 32'h00000000;
        InputData[7263:7232] = 32'h00000000;
        InputData[7295:7264] = 32'h00000000;
        InputData[7327:7296] = 32'h00000000;
        InputData[7359:7328] = 32'h00000000;
        InputData[7391:7360] = 32'h00000000;
        InputData[7423:7392] = 32'h00000000;
        InputData[7455:7424] = 32'h00000000;
        InputData[7487:7456] = 32'h00000000;
        InputData[7519:7488] = 32'h00000000;
        InputData[7551:7520] = 32'h3f800000;
        InputData[7583:7552] = 32'h3f800000;
        InputData[7615:7584] = 32'h3f800000;
        InputData[7647:7616] = 32'h00000000;
        InputData[7679:7648] = 32'h00000000;
        InputData[7711:7680] = 32'h00000000;
        InputData[7743:7712] = 32'h00000000;
        InputData[7775:7744] = 32'h3f800000;
        InputData[7807:7776] = 32'h3f800000;
        InputData[7839:7808] = 32'h3f800000;
        InputData[7871:7840] = 32'h3f800000;
        InputData[7903:7872] = 32'h3f800000;
        InputData[7935:7904] = 32'h00000000;
        InputData[7967:7936] = 32'h00000000;
        InputData[7999:7968] = 32'h00000000;
        InputData[8031:8000] = 32'h00000000;
        InputData[8063:8032] = 32'h00000000;
        InputData[8095:8064] = 32'h00000000;
        InputData[8127:8096] = 32'h00000000;
        InputData[8159:8128] = 32'h00000000;
        InputData[8191:8160] = 32'h00000000;
        InputData[8223:8192] = 32'h00000000;
        InputData[8255:8224] = 32'h00000000;
        InputData[8287:8256] = 32'h00000000;
        InputData[8319:8288] = 32'h00000000;
        InputData[8351:8320] = 32'h00000000;
        InputData[8383:8352] = 32'h00000000;
        InputData[8415:8384] = 32'h3f800000;
        InputData[8447:8416] = 32'h3f800000;
        InputData[8479:8448] = 32'h3f800000;
        InputData[8511:8480] = 32'h3f800000;
        InputData[8543:8512] = 32'h00000000;
        InputData[8575:8544] = 32'h00000000;
        InputData[8607:8576] = 32'h00000000;
        InputData[8639:8608] = 32'h3f800000;
        InputData[8671:8640] = 32'h3f800000;
        InputData[8703:8672] = 32'h3f800000;
        InputData[8735:8704] = 32'h3f800000;
        InputData[8767:8736] = 32'h3f800000;
        InputData[8799:8768] = 32'h00000000;
        InputData[8831:8800] = 32'h00000000;
        InputData[8863:8832] = 32'h00000000;
        InputData[8895:8864] = 32'h00000000;
        InputData[8927:8896] = 32'h00000000;
        InputData[8959:8928] = 32'h00000000;
        InputData[8991:8960] = 32'h00000000;
        InputData[9023:8992] = 32'h00000000;
        InputData[9055:9024] = 32'h00000000;
        InputData[9087:9056] = 32'h00000000;
        InputData[9119:9088] = 32'h00000000;
        InputData[9151:9120] = 32'h00000000;
        InputData[9183:9152] = 32'h00000000;
        InputData[9215:9184] = 32'h00000000;
        InputData[9247:9216] = 32'h00000000;
        InputData[9279:9248] = 32'h00000000;
        InputData[9311:9280] = 32'h3f800000;
        InputData[9343:9312] = 32'h3f800000;
        InputData[9375:9344] = 32'h3f800000;
        InputData[9407:9376] = 32'h00000000;
        InputData[9439:9408] = 32'h00000000;
        InputData[9471:9440] = 32'h00000000;
        InputData[9503:9472] = 32'h3f800000;
        InputData[9535:9504] = 32'h3f800000;
        InputData[9567:9536] = 32'h3f800000;
        InputData[9599:9568] = 32'h3f800000;
        InputData[9631:9600] = 32'h3f800000;
        InputData[9663:9632] = 32'h00000000;
        InputData[9695:9664] = 32'h00000000;
        InputData[9727:9696] = 32'h00000000;
        InputData[9759:9728] = 32'h00000000;
        InputData[9791:9760] = 32'h00000000;
        InputData[9823:9792] = 32'h00000000;
        InputData[9855:9824] = 32'h00000000;
        InputData[9887:9856] = 32'h00000000;
        InputData[9919:9888] = 32'h00000000;
        InputData[9951:9920] = 32'h00000000;
        InputData[9983:9952] = 32'h00000000;
        InputData[10015:9984] = 32'h00000000;
        InputData[10047:10016] = 32'h00000000;
        InputData[10079:10048] = 32'h00000000;
        InputData[10111:10080] = 32'h00000000;
        InputData[10143:10112] = 32'h00000000;
        InputData[10175:10144] = 32'h3f800000;
        InputData[10207:10176] = 32'h3f800000;
        InputData[10239:10208] = 32'h3f800000;
        InputData[10271:10240] = 32'h3f800000;
        InputData[10303:10272] = 32'h00000000;
        InputData[10335:10304] = 32'h00000000;
        InputData[10367:10336] = 32'h3f800000;
        InputData[10399:10368] = 32'h3f800000;
        InputData[10431:10400] = 32'h3f800000;
        InputData[10463:10432] = 32'h3f800000;
        InputData[10495:10464] = 32'h3f800000;
        InputData[10527:10496] = 32'h00000000;
        InputData[10559:10528] = 32'h00000000;
        InputData[10591:10560] = 32'h00000000;
        InputData[10623:10592] = 32'h00000000;
        InputData[10655:10624] = 32'h00000000;
        InputData[10687:10656] = 32'h00000000;
        InputData[10719:10688] = 32'h00000000;
        InputData[10751:10720] = 32'h00000000;
        InputData[10783:10752] = 32'h00000000;
        InputData[10815:10784] = 32'h00000000;
        InputData[10847:10816] = 32'h00000000;
        InputData[10879:10848] = 32'h00000000;
        InputData[10911:10880] = 32'h00000000;
        InputData[10943:10912] = 32'h00000000;
        InputData[10975:10944] = 32'h00000000;
        InputData[11007:10976] = 32'h00000000;
        InputData[11039:11008] = 32'h00000000;
        InputData[11071:11040] = 32'h3f800000;
        InputData[11103:11072] = 32'h3f800000;
        InputData[11135:11104] = 32'h3f800000;
        InputData[11167:11136] = 32'h00000000;
        InputData[11199:11168] = 32'h3f800000;
        InputData[11231:11200] = 32'h3f800000;
        InputData[11263:11232] = 32'h3f800000;
        InputData[11295:11264] = 32'h3f800000;
        InputData[11327:11296] = 32'h3f800000;
        InputData[11359:11328] = 32'h3f800000;
        InputData[11391:11360] = 32'h00000000;
        InputData[11423:11392] = 32'h00000000;
        InputData[11455:11424] = 32'h00000000;
        InputData[11487:11456] = 32'h00000000;
        InputData[11519:11488] = 32'h00000000;
        InputData[11551:11520] = 32'h00000000;
        InputData[11583:11552] = 32'h00000000;
        InputData[11615:11584] = 32'h00000000;
        InputData[11647:11616] = 32'h00000000;
        InputData[11679:11648] = 32'h00000000;
        InputData[11711:11680] = 32'h00000000;
        InputData[11743:11712] = 32'h00000000;
        InputData[11775:11744] = 32'h00000000;
        InputData[11807:11776] = 32'h00000000;
        InputData[11839:11808] = 32'h00000000;
        InputData[11871:11840] = 32'h00000000;
        InputData[11903:11872] = 32'h00000000;
        InputData[11935:11904] = 32'h00000000;
        InputData[11967:11936] = 32'h3f800000;
        InputData[11999:11968] = 32'h3f800000;
        InputData[12031:12000] = 32'h3f800000;
        InputData[12063:12032] = 32'h3f800000;
        InputData[12095:12064] = 32'h3f800000;
        InputData[12127:12096] = 32'h3f800000;
        InputData[12159:12128] = 32'h3f800000;
        InputData[12191:12160] = 32'h3f800000;
        InputData[12223:12192] = 32'h3f800000;
        InputData[12255:12224] = 32'h00000000;
        InputData[12287:12256] = 32'h00000000;
        InputData[12319:12288] = 32'h00000000;
        InputData[12351:12320] = 32'h00000000;
        InputData[12383:12352] = 32'h00000000;
        InputData[12415:12384] = 32'h00000000;
        InputData[12447:12416] = 32'h00000000;
        InputData[12479:12448] = 32'h00000000;
        InputData[12511:12480] = 32'h00000000;
        InputData[12543:12512] = 32'h00000000;
        InputData[12575:12544] = 32'h00000000;
        InputData[12607:12576] = 32'h00000000;
        InputData[12639:12608] = 32'h00000000;
        InputData[12671:12640] = 32'h00000000;
        InputData[12703:12672] = 32'h00000000;
        InputData[12735:12704] = 32'h00000000;
        InputData[12767:12736] = 32'h00000000;
        InputData[12799:12768] = 32'h00000000;
        InputData[12831:12800] = 32'h3f800000;
        InputData[12863:12832] = 32'h3f800000;
        InputData[12895:12864] = 32'h3f800000;
        InputData[12927:12896] = 32'h3f800000;
        InputData[12959:12928] = 32'h3f800000;
        InputData[12991:12960] = 32'h3f800000;
        InputData[13023:12992] = 32'h3f800000;
        InputData[13055:13024] = 32'h3f800000;
        InputData[13087:13056] = 32'h00000000;
        InputData[13119:13088] = 32'h00000000;
        InputData[13151:13120] = 32'h00000000;
        InputData[13183:13152] = 32'h00000000;
        InputData[13215:13184] = 32'h00000000;
        InputData[13247:13216] = 32'h00000000;
        InputData[13279:13248] = 32'h00000000;
        InputData[13311:13280] = 32'h00000000;
        InputData[13343:13312] = 32'h00000000;
        InputData[13375:13344] = 32'h00000000;
        InputData[13407:13376] = 32'h00000000;
        InputData[13439:13408] = 32'h00000000;
        InputData[13471:13440] = 32'h00000000;
        InputData[13503:13472] = 32'h00000000;
        InputData[13535:13504] = 32'h00000000;
        InputData[13567:13536] = 32'h00000000;
        InputData[13599:13568] = 32'h00000000;
        InputData[13631:13600] = 32'h00000000;
        InputData[13663:13632] = 32'h00000000;
        InputData[13695:13664] = 32'h00000000;
        InputData[13727:13696] = 32'h3f800000;
        InputData[13759:13728] = 32'h3f800000;
        InputData[13791:13760] = 32'h3f800000;
        InputData[13823:13792] = 32'h3f800000;
        InputData[13855:13824] = 32'h3f800000;
        InputData[13887:13856] = 32'h3f800000;
        InputData[13919:13888] = 32'h3f800000;
        InputData[13951:13920] = 32'h00000000;
        InputData[13983:13952] = 32'h00000000;
        InputData[14015:13984] = 32'h00000000;
        InputData[14047:14016] = 32'h00000000;
        InputData[14079:14048] = 32'h00000000;
        InputData[14111:14080] = 32'h00000000;
        InputData[14143:14112] = 32'h00000000;
        InputData[14175:14144] = 32'h00000000;
        InputData[14207:14176] = 32'h00000000;
        InputData[14239:14208] = 32'h00000000;
        InputData[14271:14240] = 32'h00000000;
        InputData[14303:14272] = 32'h00000000;
        InputData[14335:14304] = 32'h00000000;
        InputData[14367:14336] = 32'h00000000;
        InputData[14399:14368] = 32'h00000000;
        InputData[14431:14400] = 32'h00000000;
        InputData[14463:14432] = 32'h00000000;
        InputData[14495:14464] = 32'h00000000;
        InputData[14527:14496] = 32'h00000000;
        InputData[14559:14528] = 32'h00000000;
        InputData[14591:14560] = 32'h3f800000;
        InputData[14623:14592] = 32'h3f800000;
        InputData[14655:14624] = 32'h3f800000;
        InputData[14687:14656] = 32'h3f800000;
        InputData[14719:14688] = 32'h3f800000;
        InputData[14751:14720] = 32'h3f800000;
        InputData[14783:14752] = 32'h3f800000;
        InputData[14815:14784] = 32'h3f800000;
        InputData[14847:14816] = 32'h00000000;
        InputData[14879:14848] = 32'h00000000;
        InputData[14911:14880] = 32'h00000000;
        InputData[14943:14912] = 32'h00000000;
        InputData[14975:14944] = 32'h00000000;
        InputData[15007:14976] = 32'h00000000;
        InputData[15039:15008] = 32'h00000000;
        InputData[15071:15040] = 32'h00000000;
        InputData[15103:15072] = 32'h00000000;
        InputData[15135:15104] = 32'h00000000;
        InputData[15167:15136] = 32'h00000000;
        InputData[15199:15168] = 32'h00000000;
        InputData[15231:15200] = 32'h00000000;
        InputData[15263:15232] = 32'h00000000;
        InputData[15295:15264] = 32'h00000000;
        InputData[15327:15296] = 32'h00000000;
        InputData[15359:15328] = 32'h00000000;
        InputData[15391:15360] = 32'h00000000;
        InputData[15423:15392] = 32'h00000000;
        InputData[15455:15424] = 32'h00000000;
        InputData[15487:15456] = 32'h3f800000;
        InputData[15519:15488] = 32'h3f800000;
        InputData[15551:15520] = 32'h3f800000;
        InputData[15583:15552] = 32'h00000000;
        InputData[15615:15584] = 32'h3f800000;
        InputData[15647:15616] = 32'h3f800000;
        InputData[15679:15648] = 32'h3f800000;
        InputData[15711:15680] = 32'h3f800000;
        InputData[15743:15712] = 32'h3f800000;
        InputData[15775:15744] = 32'h00000000;
        InputData[15807:15776] = 32'h00000000;
        InputData[15839:15808] = 32'h00000000;
        InputData[15871:15840] = 32'h00000000;
        InputData[15903:15872] = 32'h00000000;
        InputData[15935:15904] = 32'h00000000;
        InputData[15967:15936] = 32'h00000000;
        InputData[15999:15968] = 32'h00000000;
        InputData[16031:16000] = 32'h00000000;
        InputData[16063:16032] = 32'h00000000;
        InputData[16095:16064] = 32'h00000000;
        InputData[16127:16096] = 32'h00000000;
        InputData[16159:16128] = 32'h00000000;
        InputData[16191:16160] = 32'h00000000;
        InputData[16223:16192] = 32'h00000000;
        InputData[16255:16224] = 32'h00000000;
        InputData[16287:16256] = 32'h00000000;
        InputData[16319:16288] = 32'h00000000;
        InputData[16351:16320] = 32'h3f800000;
        InputData[16383:16352] = 32'h3f800000;
        InputData[16415:16384] = 32'h3f800000;
        InputData[16447:16416] = 32'h3f800000;
        InputData[16479:16448] = 32'h00000000;
        InputData[16511:16480] = 32'h00000000;
        InputData[16543:16512] = 32'h3f800000;
        InputData[16575:16544] = 32'h3f800000;
        InputData[16607:16576] = 32'h3f800000;
        InputData[16639:16608] = 32'h3f800000;
        InputData[16671:16640] = 32'h3f800000;
        InputData[16703:16672] = 32'h00000000;
        InputData[16735:16704] = 32'h00000000;
        InputData[16767:16736] = 32'h00000000;
        InputData[16799:16768] = 32'h00000000;
        InputData[16831:16800] = 32'h00000000;
        InputData[16863:16832] = 32'h00000000;
        InputData[16895:16864] = 32'h00000000;
        InputData[16927:16896] = 32'h00000000;
        InputData[16959:16928] = 32'h00000000;
        InputData[16991:16960] = 32'h00000000;
        InputData[17023:16992] = 32'h00000000;
        InputData[17055:17024] = 32'h00000000;
        InputData[17087:17056] = 32'h00000000;
        InputData[17119:17088] = 32'h00000000;
        InputData[17151:17120] = 32'h00000000;
        InputData[17183:17152] = 32'h00000000;
        InputData[17215:17184] = 32'h00000000;
        InputData[17247:17216] = 32'h3f800000;
        InputData[17279:17248] = 32'h3f800000;
        InputData[17311:17280] = 32'h3f800000;
        InputData[17343:17312] = 32'h00000000;
        InputData[17375:17344] = 32'h00000000;
        InputData[17407:17376] = 32'h00000000;
        InputData[17439:17408] = 32'h00000000;
        InputData[17471:17440] = 32'h3f800000;
        InputData[17503:17472] = 32'h3f800000;
        InputData[17535:17504] = 32'h3f800000;
        InputData[17567:17536] = 32'h3f800000;
        InputData[17599:17568] = 32'h3f800000;
        InputData[17631:17600] = 32'h00000000;
        InputData[17663:17632] = 32'h00000000;
        InputData[17695:17664] = 32'h00000000;
        InputData[17727:17696] = 32'h00000000;
        InputData[17759:17728] = 32'h00000000;
        InputData[17791:17760] = 32'h00000000;
        InputData[17823:17792] = 32'h00000000;
        InputData[17855:17824] = 32'h00000000;
        InputData[17887:17856] = 32'h00000000;
        InputData[17919:17888] = 32'h00000000;
        InputData[17951:17920] = 32'h00000000;
        InputData[17983:17952] = 32'h00000000;
        InputData[18015:17984] = 32'h00000000;
        InputData[18047:18016] = 32'h00000000;
        InputData[18079:18048] = 32'h00000000;
        InputData[18111:18080] = 32'h3f800000;
        InputData[18143:18112] = 32'h3f800000;
        InputData[18175:18144] = 32'h3f800000;
        InputData[18207:18176] = 32'h3f800000;
        InputData[18239:18208] = 32'h00000000;
        InputData[18271:18240] = 32'h00000000;
        InputData[18303:18272] = 32'h00000000;
        InputData[18335:18304] = 32'h00000000;
        InputData[18367:18336] = 32'h00000000;
        InputData[18399:18368] = 32'h3f800000;
        InputData[18431:18400] = 32'h3f800000;
        InputData[18463:18432] = 32'h3f800000;
        InputData[18495:18464] = 32'h3f800000;
        InputData[18527:18496] = 32'h00000000;
        InputData[18559:18528] = 32'h00000000;
        InputData[18591:18560] = 32'h00000000;
        InputData[18623:18592] = 32'h00000000;
        InputData[18655:18624] = 32'h00000000;
        InputData[18687:18656] = 32'h00000000;
        InputData[18719:18688] = 32'h00000000;
        InputData[18751:18720] = 32'h00000000;
        InputData[18783:18752] = 32'h00000000;
        InputData[18815:18784] = 32'h00000000;
        InputData[18847:18816] = 32'h00000000;
        InputData[18879:18848] = 32'h00000000;
        InputData[18911:18880] = 32'h00000000;
        InputData[18943:18912] = 32'h00000000;
        InputData[18975:18944] = 32'h00000000;
        InputData[19007:18976] = 32'h3f800000;
        InputData[19039:19008] = 32'h3f800000;
        InputData[19071:19040] = 32'h3f800000;
        InputData[19103:19072] = 32'h00000000;
        InputData[19135:19104] = 32'h00000000;
        InputData[19167:19136] = 32'h00000000;
        InputData[19199:19168] = 32'h00000000;
        InputData[19231:19200] = 32'h00000000;
        InputData[19263:19232] = 32'h00000000;
        InputData[19295:19264] = 32'h00000000;
        InputData[19327:19296] = 32'h3f800000;
        InputData[19359:19328] = 32'h3f800000;
        InputData[19391:19360] = 32'h3f800000;
        InputData[19423:19392] = 32'h3f800000;
        InputData[19455:19424] = 32'h00000000;
        InputData[19487:19456] = 32'h00000000;
        InputData[19519:19488] = 32'h00000000;
        InputData[19551:19520] = 32'h00000000;
        InputData[19583:19552] = 32'h00000000;
        InputData[19615:19584] = 32'h00000000;
        InputData[19647:19616] = 32'h00000000;
        InputData[19679:19648] = 32'h00000000;
        InputData[19711:19680] = 32'h00000000;
        InputData[19743:19712] = 32'h00000000;
        InputData[19775:19744] = 32'h00000000;
        InputData[19807:19776] = 32'h00000000;
        InputData[19839:19808] = 32'h00000000;
        InputData[19871:19840] = 32'h00000000;
        InputData[19903:19872] = 32'h3f800000;
        InputData[19935:19904] = 32'h3f800000;
        InputData[19967:19936] = 32'h3f800000;
        InputData[19999:19968] = 32'h00000000;
        InputData[20031:20000] = 32'h00000000;
        InputData[20063:20032] = 32'h00000000;
        InputData[20095:20064] = 32'h00000000;
        InputData[20127:20096] = 32'h00000000;
        InputData[20159:20128] = 32'h00000000;
        InputData[20191:20160] = 32'h00000000;
        InputData[20223:20192] = 32'h00000000;
        InputData[20255:20224] = 32'h3f800000;
        InputData[20287:20256] = 32'h3f800000;
        InputData[20319:20288] = 32'h3f800000;
        InputData[20351:20320] = 32'h00000000;
        InputData[20383:20352] = 32'h00000000;
        InputData[20415:20384] = 32'h00000000;
        InputData[20447:20416] = 32'h00000000;
        InputData[20479:20448] = 32'h00000000;
        InputData[20511:20480] = 32'h00000000;
        InputData[20543:20512] = 32'h00000000;
        InputData[20575:20544] = 32'h00000000;
        InputData[20607:20576] = 32'h00000000;
        InputData[20639:20608] = 32'h00000000;
        InputData[20671:20640] = 32'h00000000;
        InputData[20703:20672] = 32'h00000000;
        InputData[20735:20704] = 32'h00000000;
        InputData[20767:20736] = 32'h00000000;
        InputData[20799:20768] = 32'h3f800000;
        InputData[20831:20800] = 32'h3f800000;
        InputData[20863:20832] = 32'h3f800000;
        InputData[20895:20864] = 32'h00000000;
        InputData[20927:20896] = 32'h00000000;
        InputData[20959:20928] = 32'h00000000;
        InputData[20991:20960] = 32'h00000000;
        InputData[21023:20992] = 32'h00000000;
        InputData[21055:21024] = 32'h00000000;
        InputData[21087:21056] = 32'h00000000;
        InputData[21119:21088] = 32'h00000000;
        InputData[21151:21120] = 32'h00000000;
        InputData[21183:21152] = 32'h3f800000;
        InputData[21215:21184] = 32'h3f800000;
        InputData[21247:21216] = 32'h00000000;
        InputData[21279:21248] = 32'h00000000;
        InputData[21311:21280] = 32'h00000000;
        InputData[21343:21312] = 32'h00000000;
        InputData[21375:21344] = 32'h00000000;
        InputData[21407:21376] = 32'h00000000;
        InputData[21439:21408] = 32'h00000000;
        InputData[21471:21440] = 32'h00000000;
        InputData[21503:21472] = 32'h00000000;
        InputData[21535:21504] = 32'h00000000;
        InputData[21567:21536] = 32'h00000000;
        InputData[21599:21568] = 32'h00000000;
        InputData[21631:21600] = 32'h00000000;
        InputData[21663:21632] = 32'h00000000;
        InputData[21695:21664] = 32'h00000000;
        InputData[21727:21696] = 32'h00000000;
        InputData[21759:21728] = 32'h00000000;
        InputData[21791:21760] = 32'h00000000;
        InputData[21823:21792] = 32'h00000000;
        InputData[21855:21824] = 32'h00000000;
        InputData[21887:21856] = 32'h00000000;
        InputData[21919:21888] = 32'h00000000;
        InputData[21951:21920] = 32'h00000000;
        InputData[21983:21952] = 32'h00000000;
        InputData[22015:21984] = 32'h00000000;
        InputData[22047:22016] = 32'h00000000;
        InputData[22079:22048] = 32'h00000000;
        InputData[22111:22080] = 32'h00000000;
        InputData[22143:22112] = 32'h00000000;
        InputData[22175:22144] = 32'h00000000;
        InputData[22207:22176] = 32'h00000000;
        InputData[22239:22208] = 32'h00000000;
        InputData[22271:22240] = 32'h00000000;
        InputData[22303:22272] = 32'h00000000;
        InputData[22335:22304] = 32'h00000000;
        InputData[22367:22336] = 32'h00000000;
        InputData[22399:22368] = 32'h00000000;
        InputData[22431:22400] = 32'h00000000;
        InputData[22463:22432] = 32'h00000000;
        InputData[22495:22464] = 32'h00000000;
        InputData[22527:22496] = 32'h00000000;
        InputData[22559:22528] = 32'h00000000;
        InputData[22591:22560] = 32'h00000000;
        InputData[22623:22592] = 32'h00000000;
        InputData[22655:22624] = 32'h00000000;
        InputData[22687:22656] = 32'h00000000;
        InputData[22719:22688] = 32'h00000000;
        InputData[22751:22720] = 32'h00000000;
        InputData[22783:22752] = 32'h00000000;
        InputData[22815:22784] = 32'h00000000;
        InputData[22847:22816] = 32'h00000000;
        InputData[22879:22848] = 32'h00000000;
        InputData[22911:22880] = 32'h00000000;
        InputData[22943:22912] = 32'h00000000;
        InputData[22975:22944] = 32'h00000000;
        InputData[23007:22976] = 32'h00000000;
        InputData[23039:23008] = 32'h00000000;
        InputData[23071:23040] = 32'h00000000;
        InputData[23103:23072] = 32'h00000000;
        InputData[23135:23104] = 32'h00000000;
        InputData[23167:23136] = 32'h00000000;
        InputData[23199:23168] = 32'h00000000;
        InputData[23231:23200] = 32'h00000000;
        InputData[23263:23232] = 32'h00000000;
        InputData[23295:23264] = 32'h00000000;
        InputData[23327:23296] = 32'h00000000;
        InputData[23359:23328] = 32'h00000000;
        InputData[23391:23360] = 32'h00000000;
        InputData[23423:23392] = 32'h00000000;
        InputData[23455:23424] = 32'h00000000;
        InputData[23487:23456] = 32'h00000000;
        InputData[23519:23488] = 32'h00000000;
        InputData[23551:23520] = 32'h00000000;
        InputData[23583:23552] = 32'h00000000;
        InputData[23615:23584] = 32'h00000000;
        InputData[23647:23616] = 32'h00000000;
        InputData[23679:23648] = 32'h00000000;
        InputData[23711:23680] = 32'h00000000;
        InputData[23743:23712] = 32'h00000000;
        InputData[23775:23744] = 32'h00000000;
        InputData[23807:23776] = 32'h00000000;
        InputData[23839:23808] = 32'h00000000;
        InputData[23871:23840] = 32'h00000000;
        InputData[23903:23872] = 32'h00000000;
        InputData[23935:23904] = 32'h00000000;
        InputData[23967:23936] = 32'h00000000;
        InputData[23999:23968] = 32'h00000000;
        InputData[24031:24000] = 32'h00000000;
        InputData[24063:24032] = 32'h00000000;
        InputData[24095:24064] = 32'h00000000;
        InputData[24127:24096] = 32'h00000000;
        InputData[24159:24128] = 32'h00000000;
        InputData[24191:24160] = 32'h00000000;
        InputData[24223:24192] = 32'h00000000;
        InputData[24255:24224] = 32'h00000000;
        InputData[24287:24256] = 32'h00000000;
        InputData[24319:24288] = 32'h00000000;
        InputData[24351:24320] = 32'h00000000;
        InputData[24383:24352] = 32'h00000000;
        InputData[24415:24384] = 32'h00000000;
        InputData[24447:24416] = 32'h00000000;
        InputData[24479:24448] = 32'h00000000;
        InputData[24511:24480] = 32'h00000000;
        InputData[24543:24512] = 32'h00000000;
        InputData[24575:24544] = 32'h00000000;
        InputData[24607:24576] = 32'h00000000;
        InputData[24639:24608] = 32'h00000000;
        InputData[24671:24640] = 32'h00000000;
        InputData[24703:24672] = 32'h00000000;
        InputData[24735:24704] = 32'h00000000;
        InputData[24767:24736] = 32'h00000000;
        InputData[24799:24768] = 32'h00000000;
        InputData[24831:24800] = 32'h00000000;
        InputData[24863:24832] = 32'h00000000;
        InputData[24895:24864] = 32'h00000000;
        InputData[24927:24896] = 32'h00000000;
        InputData[24959:24928] = 32'h00000000;
        InputData[24991:24960] = 32'h00000000;
        InputData[25023:24992] = 32'h00000000;
        InputData[25055:25024] = 32'h00000000;
        InputData[25087:25056] = 32'h00000000;
        #10000 rst = 1'b0;    
    end
    always #1 clk=~clk;
    
//    Subber ss(.X(32'hff7fffff),.Y(32'h7f7fffff),.Result(Result));
//    Adder aa(.a(32'hBFC00000),.b(32'hBFC00000),.out(Result));
//    Multiplier mm(.X(32'h1E3CE509),.Y(32'h1E3CE509),.Result(Result),.inf(inf),.overflow(overflow),.underflow(underflow));
//    Division dd(.X(32'hC115999A),.Y(32'h00000001),.Result(Result));
//    float_to_i f2i(.in(32'hff800000),.out(Result),.overflow(overflow),.underflow(underflow));
//    i_to_float i2f(.in(32'h7FFFF111),.out(Result));
//    ui_to_float ui2f(.in(32'hffff1111),.out(Result));
//    check_type ct(.in(32'hff800000),.out(Result));
    riscv_datapath_with_float riscv(.clk(clk),.rst(rst),.go(go),.frequency(2'b11),.showsel(2'b00),.IRA(1'b0),.IRB(1'b0),.IRC(1'b0),.Data(InputData),.Done(done),.Res(Res));
//    riscv_datapath riscv(.clk(clk),.rst(rst),.go(go),.frequency(2'b11),.showsel(2'b00),.IRA(1'b1),.IRB(1'b1),.IRC(1'b1),.SEG(SEG),.AN(AN),.LedData(LedData),.IR(IR)); ,.IR(IR),.FMemtoReg(FMemtoReg),.FMemWrite(FMemWrite),.ALU_Src(ALU_Src),.FRegWrite(FRegWrite),.itof(itof),.ftoi(ftoi),.RegWrite(RegWrite),.ALU_OP_2(ALU_OP_2),.AinF(AinF),.BinF(BinF),.FR1out(FR1out),.FR2out(FR2out),.FR1in(FR1in),.FR2in(FR2in),.rd(rd),.FRDin(FRDin)
//    ,.IRAin(IRAin),.IRBin(IRBin),.IRCin(IRCin),.circles(circles),.IntNo(IntNo),.clrNo(clrNo),.uret(uret),.IntAddr(IntAddr),.IntrRequest(IntrRequest) .PCout(PCout), .PCin(PCin),.Jal(Jal),.Jalr(Jalr),.BJMP(BJMP),.uret(uret),.clk_n(clk_n),.halt(halt),.R1in(R1in),.R1out(R1out),.rs1(rs1),.ecall(ecall),.LedData(LedData),.ALU_result_F(ALU_result_F)
endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/10/10 12:23:40
// Design Name: 
// Module Name: MEM_RAM_FOR_F
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module MEM_RAM_FOR_F(addr,clk,rst,str,MDin,InputData,data);
    parameter DATA_WIDTH = 32;
    parameter ADDR_WIDTH = 17;
    input [ADDR_WIDTH - 1:0] addr;
    input clk,str,rst; 
    input [25087:0] InputData;
    input [DATA_WIDTH - 1:0] MDin;
    output reg[DATA_WIDTH - 1:0] data;
    (*ram_style = "block"*) reg [DATA_WIDTH-1:0] ram[2**ADDR_WIDTH-1:0];
   
    reg [ADDR_WIDTH - 1:0] InputAddr;
    reg [25087:0] tmp;
    
    initial begin
//        begin:block_1
//            integer i;
//            for(i = 0; i < 2**ADDR_WIDTH; i = i + 1)
//            begin
//                ram[i] = 0;
//            end
//        end
//        assign InputAddr = 20'd324504;
//        assign InputAddr = 17'd81126;
        assign InputAddr = 17'd82150;
        assign tmp = InputData;
        begin: block_4
//            $readmemh("D:/CO_Team_Data/fc1_weight.hex",ram,0);//fc1_weight
//            $readmemh("D:/CO_Team_Data/fc1_bias.hex",ram,313600);//fc1_bias
//            $readmemh("D:/CO_Team_Data/fc2_weight.hex",ram,314000);//fc2_weight
//            $readmemh("D:/CO_Team_Data/fc2_bias.hex",ram,324400);//fc2_bias

//            $readmemh("D:/CO_Team_Data/fc1_weight.hex",ram,0);//fc1_weight
//            $readmemh("D:/CO_Team_Data/fc1_bias.hex",ram,78400);//fc1_bias
//            $readmemh("D:/CO_Team_Data/fc2_weight.hex",ram,78500);//fc2_weight
//            $readmemh("D:/CO_Team_Data/fc2_bias.hex",ram,81100);//fc2_bias

            $readmemh("D:/CO_Team_Data/fc1_weight.hex",ram,1024);//fc1_weight
            $readmemh("D:/CO_Team_Data/fc1_bias.hex",ram,79424);//fc1_bias
            $readmemh("D:/CO_Team_Data/fc2_weight.hex",ram,79524);//fc2_weight
            $readmemh("D:/CO_Team_Data/fc2_bias.hex",ram,82124);//
        end
    end
    
//    always@(posedge clk)
//    begin: block_3
//        ram[81126] <= InputData[31:0];
//        ram[81127] <= InputData[63:32];
//        ram[81128] <= InputData[95:64];
//        ram[81129] <= InputData[127:96];
//        ram[81130] <= InputData[159:128];
//        ram[81131] <= InputData[191:160];
//        ram[81132] <= InputData[223:192];
//        ram[81133] <= InputData[255:224];
//        ram[81134] <= InputData[287:256];
//        ram[81135] <= InputData[319:288];
//        ram[81136] <= InputData[351:320];
//        ram[81137] <= InputData[383:352];
//        ram[81138] <= InputData[415:384];
//        ram[81139] <= InputData[447:416];
//        ram[81140] <= InputData[479:448];
//        ram[81141] <= InputData[511:480];
//        ram[81142] <= InputData[543:512];
//        ram[81143] <= InputData[575:544];
//        ram[81144] <= InputData[607:576];
//        ram[81145] <= InputData[639:608];
//        ram[81146] <= InputData[671:640];
//        ram[81147] <= InputData[703:672];
//        ram[81148] <= InputData[735:704];
//        ram[81149] <= InputData[767:736];
//        ram[81150] <= InputData[799:768];
//        ram[81151] <= InputData[831:800];
//        ram[81152] <= InputData[863:832];
//        ram[81153] <= InputData[895:864];
//        ram[81154] <= InputData[927:896];
//        ram[81155] <= InputData[959:928];
//        ram[81156] <= InputData[991:960];
//        ram[81157] <= InputData[1023:992];
//        ram[81158] <= InputData[1055:1024];
//        ram[81159] <= InputData[1087:1056];
//        ram[81160] <= InputData[1119:1088];
//        ram[81161] <= InputData[1151:1120];
//        ram[81162] <= InputData[1183:1152];
//        ram[81163] <= InputData[1215:1184];
//        ram[81164] <= InputData[1247:1216];
//        ram[81165] <= InputData[1279:1248];
//        ram[81166] <= InputData[1311:1280];
//        ram[81167] <= InputData[1343:1312];
//        ram[81168] <= InputData[1375:1344];
//        ram[81169] <= InputData[1407:1376];
//        ram[81170] <= InputData[1439:1408];
//        ram[81171] <= InputData[1471:1440];
//        ram[81172] <= InputData[1503:1472];
//        ram[81173] <= InputData[1535:1504];
//        ram[81174] <= InputData[1567:1536];
//        ram[81175] <= InputData[1599:1568];
//        ram[81176] <= InputData[1631:1600];
//        ram[81177] <= InputData[1663:1632];
//        ram[81178] <= InputData[1695:1664];
//        ram[81179] <= InputData[1727:1696];
//        ram[81180] <= InputData[1759:1728];
//        ram[81181] <= InputData[1791:1760];
//        ram[81182] <= InputData[1823:1792];
//        ram[81183] <= InputData[1855:1824];
//        ram[81184] <= InputData[1887:1856];
//        ram[81185] <= InputData[1919:1888];
//        ram[81186] <= InputData[1951:1920];
//        ram[81187] <= InputData[1983:1952];
//        ram[81188] <= InputData[2015:1984];
//        ram[81189] <= InputData[2047:2016];
//        ram[81190] <= InputData[2079:2048];
//        ram[81191] <= InputData[2111:2080];
//        ram[81192] <= InputData[2143:2112];
//        ram[81193] <= InputData[2175:2144];
//        ram[81194] <= InputData[2207:2176];
//        ram[81195] <= InputData[2239:2208];
//        ram[81196] <= InputData[2271:2240];
//        ram[81197] <= InputData[2303:2272];
//        ram[81198] <= InputData[2335:2304];
//        ram[81199] <= InputData[2367:2336];
//        ram[81200] <= InputData[2399:2368];
//        ram[81201] <= InputData[2431:2400];
//        ram[81202] <= InputData[2463:2432];
//        ram[81203] <= InputData[2495:2464];
//        ram[81204] <= InputData[2527:2496];
//        ram[81205] <= InputData[2559:2528];
//        ram[81206] <= InputData[2591:2560];
//        ram[81207] <= InputData[2623:2592];
//        ram[81208] <= InputData[2655:2624];
//        ram[81209] <= InputData[2687:2656];
//        ram[81210] <= InputData[2719:2688];
//        ram[81211] <= InputData[2751:2720];
//        ram[81212] <= InputData[2783:2752];
//        ram[81213] <= InputData[2815:2784];
//        ram[81214] <= InputData[2847:2816];
//        ram[81215] <= InputData[2879:2848];
//        ram[81216] <= InputData[2911:2880];
//        ram[81217] <= InputData[2943:2912];
//        ram[81218] <= InputData[2975:2944];
//        ram[81219] <= InputData[3007:2976];
//        ram[81220] <= InputData[3039:3008];
//        ram[81221] <= InputData[3071:3040];
//        ram[81222] <= InputData[3103:3072];
//        ram[81223] <= InputData[3135:3104];
//        ram[81224] <= InputData[3167:3136];
//        ram[81225] <= InputData[3199:3168];
//        ram[81226] <= InputData[3231:3200];
//        ram[81227] <= InputData[3263:3232];
//        ram[81228] <= InputData[3295:3264];
//        ram[81229] <= InputData[3327:3296];
//        ram[81230] <= InputData[3359:3328];
//        ram[81231] <= InputData[3391:3360];
//        ram[81232] <= InputData[3423:3392];
//        ram[81233] <= InputData[3455:3424];
//        ram[81234] <= InputData[3487:3456];
//        ram[81235] <= InputData[3519:3488];
//        ram[81236] <= InputData[3551:3520];
//        ram[81237] <= InputData[3583:3552];
//        ram[81238] <= InputData[3615:3584];
//        ram[81239] <= InputData[3647:3616];
//        ram[81240] <= InputData[3679:3648];
//        ram[81241] <= InputData[3711:3680];
//        ram[81242] <= InputData[3743:3712];
//        ram[81243] <= InputData[3775:3744];
//        ram[81244] <= InputData[3807:3776];
//        ram[81245] <= InputData[3839:3808];
//        ram[81246] <= InputData[3871:3840];
//        ram[81247] <= InputData[3903:3872];
//        ram[81248] <= InputData[3935:3904];
//        ram[81249] <= InputData[3967:3936];
//        ram[81250] <= InputData[3999:3968];
//        ram[81251] <= InputData[4031:4000];
//        ram[81252] <= InputData[4063:4032];
//        ram[81253] <= InputData[4095:4064];
//        ram[81254] <= InputData[4127:4096];
//        ram[81255] <= InputData[4159:4128];
//        ram[81256] <= InputData[4191:4160];
//        ram[81257] <= InputData[4223:4192];
//        ram[81258] <= InputData[4255:4224];
//        ram[81259] <= InputData[4287:4256];
//        ram[81260] <= InputData[4319:4288];
//        ram[81261] <= InputData[4351:4320];
//        ram[81262] <= InputData[4383:4352];
//        ram[81263] <= InputData[4415:4384];
//        ram[81264] <= InputData[4447:4416];
//        ram[81265] <= InputData[4479:4448];
//        ram[81266] <= InputData[4511:4480];
//        ram[81267] <= InputData[4543:4512];
//        ram[81268] <= InputData[4575:4544];
//        ram[81269] <= InputData[4607:4576];
//        ram[81270] <= InputData[4639:4608];
//        ram[81271] <= InputData[4671:4640];
//        ram[81272] <= InputData[4703:4672];
//        ram[81273] <= InputData[4735:4704];
//        ram[81274] <= InputData[4767:4736];
//        ram[81275] <= InputData[4799:4768];
//        ram[81276] <= InputData[4831:4800];
//        ram[81277] <= InputData[4863:4832];
//        ram[81278] <= InputData[4895:4864];
//        ram[81279] <= InputData[4927:4896];
//        ram[81280] <= InputData[4959:4928];
//        ram[81281] <= InputData[4991:4960];
//        ram[81282] <= InputData[5023:4992];
//        ram[81283] <= InputData[5055:5024];
//        ram[81284] <= InputData[5087:5056];
//        ram[81285] <= InputData[5119:5088];
//        ram[81286] <= InputData[5151:5120];
//        ram[81287] <= InputData[5183:5152];
//        ram[81288] <= InputData[5215:5184];
//        ram[81289] <= InputData[5247:5216];
//        ram[81290] <= InputData[5279:5248];
//        ram[81291] <= InputData[5311:5280];
//        ram[81292] <= InputData[5343:5312];
//        ram[81293] <= InputData[5375:5344];
//        ram[81294] <= InputData[5407:5376];
//        ram[81295] <= InputData[5439:5408];
//        ram[81296] <= InputData[5471:5440];
//        ram[81297] <= InputData[5503:5472];
//        ram[81298] <= InputData[5535:5504];
//        ram[81299] <= InputData[5567:5536];
//        ram[81300] <= InputData[5599:5568];
//        ram[81301] <= InputData[5631:5600];
//        ram[81302] <= InputData[5663:5632];
//        ram[81303] <= InputData[5695:5664];
//        ram[81304] <= InputData[5727:5696];
//        ram[81305] <= InputData[5759:5728];
//        ram[81306] <= InputData[5791:5760];
//        ram[81307] <= InputData[5823:5792];
//        ram[81308] <= InputData[5855:5824];
//        ram[81309] <= InputData[5887:5856];
//        ram[81310] <= InputData[5919:5888];
//        ram[81311] <= InputData[5951:5920];
//        ram[81312] <= InputData[5983:5952];
//        ram[81313] <= InputData[6015:5984];
//        ram[81314] <= InputData[6047:6016];
//        ram[81315] <= InputData[6079:6048];
//        ram[81316] <= InputData[6111:6080];
//        ram[81317] <= InputData[6143:6112];
//        ram[81318] <= InputData[6175:6144];
//        ram[81319] <= InputData[6207:6176];
//        ram[81320] <= InputData[6239:6208];
//        ram[81321] <= InputData[6271:6240];
//        ram[81322] <= InputData[6303:6272];
//        ram[81323] <= InputData[6335:6304];
//        ram[81324] <= InputData[6367:6336];
//        ram[81325] <= InputData[6399:6368];
//        ram[81326] <= InputData[6431:6400];
//        ram[81327] <= InputData[6463:6432];
//        ram[81328] <= InputData[6495:6464];
//        ram[81329] <= InputData[6527:6496];
//        ram[81330] <= InputData[6559:6528];
//        ram[81331] <= InputData[6591:6560];
//        ram[81332] <= InputData[6623:6592];
//        ram[81333] <= InputData[6655:6624];
//        ram[81334] <= InputData[6687:6656];
//        ram[81335] <= InputData[6719:6688];
//        ram[81336] <= InputData[6751:6720];
//        ram[81337] <= InputData[6783:6752];
//        ram[81338] <= InputData[6815:6784];
//        ram[81339] <= InputData[6847:6816];
//        ram[81340] <= InputData[6879:6848];
//        ram[81341] <= InputData[6911:6880];
//        ram[81342] <= InputData[6943:6912];
//        ram[81343] <= InputData[6975:6944];
//        ram[81344] <= InputData[7007:6976];
//        ram[81345] <= InputData[7039:7008];
//        ram[81346] <= InputData[7071:7040];
//        ram[81347] <= InputData[7103:7072];
//        ram[81348] <= InputData[7135:7104];
//        ram[81349] <= InputData[7167:7136];
//        ram[81350] <= InputData[7199:7168];
//        ram[81351] <= InputData[7231:7200];
//        ram[81352] <= InputData[7263:7232];
//        ram[81353] <= InputData[7295:7264];
//        ram[81354] <= InputData[7327:7296];
//        ram[81355] <= InputData[7359:7328];
//        ram[81356] <= InputData[7391:7360];
//        ram[81357] <= InputData[7423:7392];
//        ram[81358] <= InputData[7455:7424];
//        ram[81359] <= InputData[7487:7456];
//        ram[81360] <= InputData[7519:7488];
//        ram[81361] <= InputData[7551:7520];
//        ram[81362] <= InputData[7583:7552];
//        ram[81363] <= InputData[7615:7584];
//        ram[81364] <= InputData[7647:7616];
//        ram[81365] <= InputData[7679:7648];
//        ram[81366] <= InputData[7711:7680];
//        ram[81367] <= InputData[7743:7712];
//        ram[81368] <= InputData[7775:7744];
//        ram[81369] <= InputData[7807:7776];
//        ram[81370] <= InputData[7839:7808];
//        ram[81371] <= InputData[7871:7840];
//        ram[81372] <= InputData[7903:7872];
//        ram[81373] <= InputData[7935:7904];
//        ram[81374] <= InputData[7967:7936];
//        ram[81375] <= InputData[7999:7968];
//        ram[81376] <= InputData[8031:8000];
//        ram[81377] <= InputData[8063:8032];
//        ram[81378] <= InputData[8095:8064];
//        ram[81379] <= InputData[8127:8096];
//        ram[81380] <= InputData[8159:8128];
//        ram[81381] <= InputData[8191:8160];
//        ram[81382] <= InputData[8223:8192];
//        ram[81383] <= InputData[8255:8224];
//        ram[81384] <= InputData[8287:8256];
//        ram[81385] <= InputData[8319:8288];
//        ram[81386] <= InputData[8351:8320];
//        ram[81387] <= InputData[8383:8352];
//        ram[81388] <= InputData[8415:8384];
//        ram[81389] <= InputData[8447:8416];
//        ram[81390] <= InputData[8479:8448];
//        ram[81391] <= InputData[8511:8480];
//        ram[81392] <= InputData[8543:8512];
//        ram[81393] <= InputData[8575:8544];
//        ram[81394] <= InputData[8607:8576];
//        ram[81395] <= InputData[8639:8608];
//        ram[81396] <= InputData[8671:8640];
//        ram[81397] <= InputData[8703:8672];
//        ram[81398] <= InputData[8735:8704];
//        ram[81399] <= InputData[8767:8736];
//        ram[81400] <= InputData[8799:8768];
//        ram[81401] <= InputData[8831:8800];
//        ram[81402] <= InputData[8863:8832];
//        ram[81403] <= InputData[8895:8864];
//        ram[81404] <= InputData[8927:8896];
//        ram[81405] <= InputData[8959:8928];
//        ram[81406] <= InputData[8991:8960];
//        ram[81407] <= InputData[9023:8992];
//        ram[81408] <= InputData[9055:9024];
//        ram[81409] <= InputData[9087:9056];
//        ram[81410] <= InputData[9119:9088];
//        ram[81411] <= InputData[9151:9120];
//        ram[81412] <= InputData[9183:9152];
//        ram[81413] <= InputData[9215:9184];
//        ram[81414] <= InputData[9247:9216];
//        ram[81415] <= InputData[9279:9248];
//        ram[81416] <= InputData[9311:9280];
//        ram[81417] <= InputData[9343:9312];
//        ram[81418] <= InputData[9375:9344];
//        ram[81419] <= InputData[9407:9376];
//        ram[81420] <= InputData[9439:9408];
//        ram[81421] <= InputData[9471:9440];
//        ram[81422] <= InputData[9503:9472];
//        ram[81423] <= InputData[9535:9504];
//        ram[81424] <= InputData[9567:9536];
//        ram[81425] <= InputData[9599:9568];
//        ram[81426] <= InputData[9631:9600];
//        ram[81427] <= InputData[9663:9632];
//        ram[81428] <= InputData[9695:9664];
//        ram[81429] <= InputData[9727:9696];
//        ram[81430] <= InputData[9759:9728];
//        ram[81431] <= InputData[9791:9760];
//        ram[81432] <= InputData[9823:9792];
//        ram[81433] <= InputData[9855:9824];
//        ram[81434] <= InputData[9887:9856];
//        ram[81435] <= InputData[9919:9888];
//        ram[81436] <= InputData[9951:9920];
//        ram[81437] <= InputData[9983:9952];
//        ram[81438] <= InputData[10015:9984];
//        ram[81439] <= InputData[10047:10016];
//        ram[81440] <= InputData[10079:10048];
//        ram[81441] <= InputData[10111:10080];
//        ram[81442] <= InputData[10143:10112];
//        ram[81443] <= InputData[10175:10144];
//        ram[81444] <= InputData[10207:10176];
//        ram[81445] <= InputData[10239:10208];
//        ram[81446] <= InputData[10271:10240];
//        ram[81447] <= InputData[10303:10272];
//        ram[81448] <= InputData[10335:10304];
//        ram[81449] <= InputData[10367:10336];
//        ram[81450] <= InputData[10399:10368];
//        ram[81451] <= InputData[10431:10400];
//        ram[81452] <= InputData[10463:10432];
//        ram[81453] <= InputData[10495:10464];
//        ram[81454] <= InputData[10527:10496];
//        ram[81455] <= InputData[10559:10528];
//        ram[81456] <= InputData[10591:10560];
//        ram[81457] <= InputData[10623:10592];
//        ram[81458] <= InputData[10655:10624];
//        ram[81459] <= InputData[10687:10656];
//        ram[81460] <= InputData[10719:10688];
//        ram[81461] <= InputData[10751:10720];
//        ram[81462] <= InputData[10783:10752];
//        ram[81463] <= InputData[10815:10784];
//        ram[81464] <= InputData[10847:10816];
//        ram[81465] <= InputData[10879:10848];
//        ram[81466] <= InputData[10911:10880];
//        ram[81467] <= InputData[10943:10912];
//        ram[81468] <= InputData[10975:10944];
//        ram[81469] <= InputData[11007:10976];
//        ram[81470] <= InputData[11039:11008];
//        ram[81471] <= InputData[11071:11040];
//        ram[81472] <= InputData[11103:11072];
//        ram[81473] <= InputData[11135:11104];
//        ram[81474] <= InputData[11167:11136];
//        ram[81475] <= InputData[11199:11168];
//        ram[81476] <= InputData[11231:11200];
//        ram[81477] <= InputData[11263:11232];
//        ram[81478] <= InputData[11295:11264];
//        ram[81479] <= InputData[11327:11296];
//        ram[81480] <= InputData[11359:11328];
//        ram[81481] <= InputData[11391:11360];
//        ram[81482] <= InputData[11423:11392];
//        ram[81483] <= InputData[11455:11424];
//        ram[81484] <= InputData[11487:11456];
//        ram[81485] <= InputData[11519:11488];
//        ram[81486] <= InputData[11551:11520];
//        ram[81487] <= InputData[11583:11552];
//        ram[81488] <= InputData[11615:11584];
//        ram[81489] <= InputData[11647:11616];
//        ram[81490] <= InputData[11679:11648];
//        ram[81491] <= InputData[11711:11680];
//        ram[81492] <= InputData[11743:11712];
//        ram[81493] <= InputData[11775:11744];
//        ram[81494] <= InputData[11807:11776];
//        ram[81495] <= InputData[11839:11808];
//        ram[81496] <= InputData[11871:11840];
//        ram[81497] <= InputData[11903:11872];
//        ram[81498] <= InputData[11935:11904];
//        ram[81499] <= InputData[11967:11936];
//        ram[81500] <= InputData[11999:11968];
//        ram[81501] <= InputData[12031:12000];
//        ram[81502] <= InputData[12063:12032];
//        ram[81503] <= InputData[12095:12064];
//        ram[81504] <= InputData[12127:12096];
//        ram[81505] <= InputData[12159:12128];
//        ram[81506] <= InputData[12191:12160];
//        ram[81507] <= InputData[12223:12192];
//        ram[81508] <= InputData[12255:12224];
//        ram[81509] <= InputData[12287:12256];
//        ram[81510] <= InputData[12319:12288];
//        ram[81511] <= InputData[12351:12320];
//        ram[81512] <= InputData[12383:12352];
//        ram[81513] <= InputData[12415:12384];
//        ram[81514] <= InputData[12447:12416];
//        ram[81515] <= InputData[12479:12448];
//        ram[81516] <= InputData[12511:12480];
//        ram[81517] <= InputData[12543:12512];
//        ram[81518] <= InputData[12575:12544];
//        ram[81519] <= InputData[12607:12576];
//        ram[81520] <= InputData[12639:12608];
//        ram[81521] <= InputData[12671:12640];
//        ram[81522] <= InputData[12703:12672];
//        ram[81523] <= InputData[12735:12704];
//        ram[81524] <= InputData[12767:12736];
//        ram[81525] <= InputData[12799:12768];
//        ram[81526] <= InputData[12831:12800];
//        ram[81527] <= InputData[12863:12832];
//        ram[81528] <= InputData[12895:12864];
//        ram[81529] <= InputData[12927:12896];
//        ram[81530] <= InputData[12959:12928];
//        ram[81531] <= InputData[12991:12960];
//        ram[81532] <= InputData[13023:12992];
//        ram[81533] <= InputData[13055:13024];
//        ram[81534] <= InputData[13087:13056];
//        ram[81535] <= InputData[13119:13088];
//        ram[81536] <= InputData[13151:13120];
//        ram[81537] <= InputData[13183:13152];
//        ram[81538] <= InputData[13215:13184];
//        ram[81539] <= InputData[13247:13216];
//        ram[81540] <= InputData[13279:13248];
//        ram[81541] <= InputData[13311:13280];
//        ram[81542] <= InputData[13343:13312];
//        ram[81543] <= InputData[13375:13344];
//        ram[81544] <= InputData[13407:13376];
//        ram[81545] <= InputData[13439:13408];
//        ram[81546] <= InputData[13471:13440];
//        ram[81547] <= InputData[13503:13472];
//        ram[81548] <= InputData[13535:13504];
//        ram[81549] <= InputData[13567:13536];
//        ram[81550] <= InputData[13599:13568];
//        ram[81551] <= InputData[13631:13600];
//        ram[81552] <= InputData[13663:13632];
//        ram[81553] <= InputData[13695:13664];
//        ram[81554] <= InputData[13727:13696];
//        ram[81555] <= InputData[13759:13728];
//        ram[81556] <= InputData[13791:13760];
//        ram[81557] <= InputData[13823:13792];
//        ram[81558] <= InputData[13855:13824];
//        ram[81559] <= InputData[13887:13856];
//        ram[81560] <= InputData[13919:13888];
//        ram[81561] <= InputData[13951:13920];
//        ram[81562] <= InputData[13983:13952];
//        ram[81563] <= InputData[14015:13984];
//        ram[81564] <= InputData[14047:14016];
//        ram[81565] <= InputData[14079:14048];
//        ram[81566] <= InputData[14111:14080];
//        ram[81567] <= InputData[14143:14112];
//        ram[81568] <= InputData[14175:14144];
//        ram[81569] <= InputData[14207:14176];
//        ram[81570] <= InputData[14239:14208];
//        ram[81571] <= InputData[14271:14240];
//        ram[81572] <= InputData[14303:14272];
//        ram[81573] <= InputData[14335:14304];
//        ram[81574] <= InputData[14367:14336];
//        ram[81575] <= InputData[14399:14368];
//        ram[81576] <= InputData[14431:14400];
//        ram[81577] <= InputData[14463:14432];
//        ram[81578] <= InputData[14495:14464];
//        ram[81579] <= InputData[14527:14496];
//        ram[81580] <= InputData[14559:14528];
//        ram[81581] <= InputData[14591:14560];
//        ram[81582] <= InputData[14623:14592];
//        ram[81583] <= InputData[14655:14624];
//        ram[81584] <= InputData[14687:14656];
//        ram[81585] <= InputData[14719:14688];
//        ram[81586] <= InputData[14751:14720];
//        ram[81587] <= InputData[14783:14752];
//        ram[81588] <= InputData[14815:14784];
//        ram[81589] <= InputData[14847:14816];
//        ram[81590] <= InputData[14879:14848];
//        ram[81591] <= InputData[14911:14880];
//        ram[81592] <= InputData[14943:14912];
//        ram[81593] <= InputData[14975:14944];
//        ram[81594] <= InputData[15007:14976];
//        ram[81595] <= InputData[15039:15008];
//        ram[81596] <= InputData[15071:15040];
//        ram[81597] <= InputData[15103:15072];
//        ram[81598] <= InputData[15135:15104];
//        ram[81599] <= InputData[15167:15136];
//        ram[81600] <= InputData[15199:15168];
//        ram[81601] <= InputData[15231:15200];
//        ram[81602] <= InputData[15263:15232];
//        ram[81603] <= InputData[15295:15264];
//        ram[81604] <= InputData[15327:15296];
//        ram[81605] <= InputData[15359:15328];
//        ram[81606] <= InputData[15391:15360];
//        ram[81607] <= InputData[15423:15392];
//        ram[81608] <= InputData[15455:15424];
//        ram[81609] <= InputData[15487:15456];
//        ram[81610] <= InputData[15519:15488];
//        ram[81611] <= InputData[15551:15520];
//        ram[81612] <= InputData[15583:15552];
//        ram[81613] <= InputData[15615:15584];
//        ram[81614] <= InputData[15647:15616];
//        ram[81615] <= InputData[15679:15648];
//        ram[81616] <= InputData[15711:15680];
//        ram[81617] <= InputData[15743:15712];
//        ram[81618] <= InputData[15775:15744];
//        ram[81619] <= InputData[15807:15776];
//        ram[81620] <= InputData[15839:15808];
//        ram[81621] <= InputData[15871:15840];
//        ram[81622] <= InputData[15903:15872];
//        ram[81623] <= InputData[15935:15904];
//        ram[81624] <= InputData[15967:15936];
//        ram[81625] <= InputData[15999:15968];
//        ram[81626] <= InputData[16031:16000];
//        ram[81627] <= InputData[16063:16032];
//        ram[81628] <= InputData[16095:16064];
//        ram[81629] <= InputData[16127:16096];
//        ram[81630] <= InputData[16159:16128];
//        ram[81631] <= InputData[16191:16160];
//        ram[81632] <= InputData[16223:16192];
//        ram[81633] <= InputData[16255:16224];
//        ram[81634] <= InputData[16287:16256];
//        ram[81635] <= InputData[16319:16288];
//        ram[81636] <= InputData[16351:16320];
//        ram[81637] <= InputData[16383:16352];
//        ram[81638] <= InputData[16415:16384];
//        ram[81639] <= InputData[16447:16416];
//        ram[81640] <= InputData[16479:16448];
//        ram[81641] <= InputData[16511:16480];
//        ram[81642] <= InputData[16543:16512];
//        ram[81643] <= InputData[16575:16544];
//        ram[81644] <= InputData[16607:16576];
//        ram[81645] <= InputData[16639:16608];
//        ram[81646] <= InputData[16671:16640];
//        ram[81647] <= InputData[16703:16672];
//        ram[81648] <= InputData[16735:16704];
//        ram[81649] <= InputData[16767:16736];
//        ram[81650] <= InputData[16799:16768];
//        ram[81651] <= InputData[16831:16800];
//        ram[81652] <= InputData[16863:16832];
//        ram[81653] <= InputData[16895:16864];
//        ram[81654] <= InputData[16927:16896];
//        ram[81655] <= InputData[16959:16928];
//        ram[81656] <= InputData[16991:16960];
//        ram[81657] <= InputData[17023:16992];
//        ram[81658] <= InputData[17055:17024];
//        ram[81659] <= InputData[17087:17056];
//        ram[81660] <= InputData[17119:17088];
//        ram[81661] <= InputData[17151:17120];
//        ram[81662] <= InputData[17183:17152];
//        ram[81663] <= InputData[17215:17184];
//        ram[81664] <= InputData[17247:17216];
//        ram[81665] <= InputData[17279:17248];
//        ram[81666] <= InputData[17311:17280];
//        ram[81667] <= InputData[17343:17312];
//        ram[81668] <= InputData[17375:17344];
//        ram[81669] <= InputData[17407:17376];
//        ram[81670] <= InputData[17439:17408];
//        ram[81671] <= InputData[17471:17440];
//        ram[81672] <= InputData[17503:17472];
//        ram[81673] <= InputData[17535:17504];
//        ram[81674] <= InputData[17567:17536];
//        ram[81675] <= InputData[17599:17568];
//        ram[81676] <= InputData[17631:17600];
//        ram[81677] <= InputData[17663:17632];
//        ram[81678] <= InputData[17695:17664];
//        ram[81679] <= InputData[17727:17696];
//        ram[81680] <= InputData[17759:17728];
//        ram[81681] <= InputData[17791:17760];
//        ram[81682] <= InputData[17823:17792];
//        ram[81683] <= InputData[17855:17824];
//        ram[81684] <= InputData[17887:17856];
//        ram[81685] <= InputData[17919:17888];
//        ram[81686] <= InputData[17951:17920];
//        ram[81687] <= InputData[17983:17952];
//        ram[81688] <= InputData[18015:17984];
//        ram[81689] <= InputData[18047:18016];
//        ram[81690] <= InputData[18079:18048];
//        ram[81691] <= InputData[18111:18080];
//        ram[81692] <= InputData[18143:18112];
//        ram[81693] <= InputData[18175:18144];
//        ram[81694] <= InputData[18207:18176];
//        ram[81695] <= InputData[18239:18208];
//        ram[81696] <= InputData[18271:18240];
//        ram[81697] <= InputData[18303:18272];
//        ram[81698] <= InputData[18335:18304];
//        ram[81699] <= InputData[18367:18336];
//        ram[81700] <= InputData[18399:18368];
//        ram[81701] <= InputData[18431:18400];
//        ram[81702] <= InputData[18463:18432];
//        ram[81703] <= InputData[18495:18464];
//        ram[81704] <= InputData[18527:18496];
//        ram[81705] <= InputData[18559:18528];
//        ram[81706] <= InputData[18591:18560];
//        ram[81707] <= InputData[18623:18592];
//        ram[81708] <= InputData[18655:18624];
//        ram[81709] <= InputData[18687:18656];
//        ram[81710] <= InputData[18719:18688];
//        ram[81711] <= InputData[18751:18720];
//        ram[81712] <= InputData[18783:18752];
//        ram[81713] <= InputData[18815:18784];
//        ram[81714] <= InputData[18847:18816];
//        ram[81715] <= InputData[18879:18848];
//        ram[81716] <= InputData[18911:18880];
//        ram[81717] <= InputData[18943:18912];
//        ram[81718] <= InputData[18975:18944];
//        ram[81719] <= InputData[19007:18976];
//        ram[81720] <= InputData[19039:19008];
//        ram[81721] <= InputData[19071:19040];
//        ram[81722] <= InputData[19103:19072];
//        ram[81723] <= InputData[19135:19104];
//        ram[81724] <= InputData[19167:19136];
//        ram[81725] <= InputData[19199:19168];
//        ram[81726] <= InputData[19231:19200];
//        ram[81727] <= InputData[19263:19232];
//        ram[81728] <= InputData[19295:19264];
//        ram[81729] <= InputData[19327:19296];
//        ram[81730] <= InputData[19359:19328];
//        ram[81731] <= InputData[19391:19360];
//        ram[81732] <= InputData[19423:19392];
//        ram[81733] <= InputData[19455:19424];
//        ram[81734] <= InputData[19487:19456];
//        ram[81735] <= InputData[19519:19488];
//        ram[81736] <= InputData[19551:19520];
//        ram[81737] <= InputData[19583:19552];
//        ram[81738] <= InputData[19615:19584];
//        ram[81739] <= InputData[19647:19616];
//        ram[81740] <= InputData[19679:19648];
//        ram[81741] <= InputData[19711:19680];
//        ram[81742] <= InputData[19743:19712];
//        ram[81743] <= InputData[19775:19744];
//        ram[81744] <= InputData[19807:19776];
//        ram[81745] <= InputData[19839:19808];
//        ram[81746] <= InputData[19871:19840];
//        ram[81747] <= InputData[19903:19872];
//        ram[81748] <= InputData[19935:19904];
//        ram[81749] <= InputData[19967:19936];
//        ram[81750] <= InputData[19999:19968];
//        ram[81751] <= InputData[20031:20000];
//        ram[81752] <= InputData[20063:20032];
//        ram[81753] <= InputData[20095:20064];
//        ram[81754] <= InputData[20127:20096];
//        ram[81755] <= InputData[20159:20128];
//        ram[81756] <= InputData[20191:20160];
//        ram[81757] <= InputData[20223:20192];
//        ram[81758] <= InputData[20255:20224];
//        ram[81759] <= InputData[20287:20256];
//        ram[81760] <= InputData[20319:20288];
//        ram[81761] <= InputData[20351:20320];
//        ram[81762] <= InputData[20383:20352];
//        ram[81763] <= InputData[20415:20384];
//        ram[81764] <= InputData[20447:20416];
//        ram[81765] <= InputData[20479:20448];
//        ram[81766] <= InputData[20511:20480];
//        ram[81767] <= InputData[20543:20512];
//        ram[81768] <= InputData[20575:20544];
//        ram[81769] <= InputData[20607:20576];
//        ram[81770] <= InputData[20639:20608];
//        ram[81771] <= InputData[20671:20640];
//        ram[81772] <= InputData[20703:20672];
//        ram[81773] <= InputData[20735:20704];
//        ram[81774] <= InputData[20767:20736];
//        ram[81775] <= InputData[20799:20768];
//        ram[81776] <= InputData[20831:20800];
//        ram[81777] <= InputData[20863:20832];
//        ram[81778] <= InputData[20895:20864];
//        ram[81779] <= InputData[20927:20896];
//        ram[81780] <= InputData[20959:20928];
//        ram[81781] <= InputData[20991:20960];
//        ram[81782] <= InputData[21023:20992];
//        ram[81783] <= InputData[21055:21024];
//        ram[81784] <= InputData[21087:21056];
//        ram[81785] <= InputData[21119:21088];
//        ram[81786] <= InputData[21151:21120];
//        ram[81787] <= InputData[21183:21152];
//        ram[81788] <= InputData[21215:21184];
//        ram[81789] <= InputData[21247:21216];
//        ram[81790] <= InputData[21279:21248];
//        ram[81791] <= InputData[21311:21280];
//        ram[81792] <= InputData[21343:21312];
//        ram[81793] <= InputData[21375:21344];
//        ram[81794] <= InputData[21407:21376];
//        ram[81795] <= InputData[21439:21408];
//        ram[81796] <= InputData[21471:21440];
//        ram[81797] <= InputData[21503:21472];
//        ram[81798] <= InputData[21535:21504];
//        ram[81799] <= InputData[21567:21536];
//        ram[81800] <= InputData[21599:21568];
//        ram[81801] <= InputData[21631:21600];
//        ram[81802] <= InputData[21663:21632];
//        ram[81803] <= InputData[21695:21664];
//        ram[81804] <= InputData[21727:21696];
//        ram[81805] <= InputData[21759:21728];
//        ram[81806] <= InputData[21791:21760];
//        ram[81807] <= InputData[21823:21792];
//        ram[81808] <= InputData[21855:21824];
//        ram[81809] <= InputData[21887:21856];
//        ram[81810] <= InputData[21919:21888];
//        ram[81811] <= InputData[21951:21920];
//        ram[81812] <= InputData[21983:21952];
//        ram[81813] <= InputData[22015:21984];
//        ram[81814] <= InputData[22047:22016];
//        ram[81815] <= InputData[22079:22048];
//        ram[81816] <= InputData[22111:22080];
//        ram[81817] <= InputData[22143:22112];
//        ram[81818] <= InputData[22175:22144];
//        ram[81819] <= InputData[22207:22176];
//        ram[81820] <= InputData[22239:22208];
//        ram[81821] <= InputData[22271:22240];
//        ram[81822] <= InputData[22303:22272];
//        ram[81823] <= InputData[22335:22304];
//        ram[81824] <= InputData[22367:22336];
//        ram[81825] <= InputData[22399:22368];
//        ram[81826] <= InputData[22431:22400];
//        ram[81827] <= InputData[22463:22432];
//        ram[81828] <= InputData[22495:22464];
//        ram[81829] <= InputData[22527:22496];
//        ram[81830] <= InputData[22559:22528];
//        ram[81831] <= InputData[22591:22560];
//        ram[81832] <= InputData[22623:22592];
//        ram[81833] <= InputData[22655:22624];
//        ram[81834] <= InputData[22687:22656];
//        ram[81835] <= InputData[22719:22688];
//        ram[81836] <= InputData[22751:22720];
//        ram[81837] <= InputData[22783:22752];
//        ram[81838] <= InputData[22815:22784];
//        ram[81839] <= InputData[22847:22816];
//        ram[81840] <= InputData[22879:22848];
//        ram[81841] <= InputData[22911:22880];
//        ram[81842] <= InputData[22943:22912];
//        ram[81843] <= InputData[22975:22944];
//        ram[81844] <= InputData[23007:22976];
//        ram[81845] <= InputData[23039:23008];
//        ram[81846] <= InputData[23071:23040];
//        ram[81847] <= InputData[23103:23072];
//        ram[81848] <= InputData[23135:23104];
//        ram[81849] <= InputData[23167:23136];
//        ram[81850] <= InputData[23199:23168];
//        ram[81851] <= InputData[23231:23200];
//        ram[81852] <= InputData[23263:23232];
//        ram[81853] <= InputData[23295:23264];
//        ram[81854] <= InputData[23327:23296];
//        ram[81855] <= InputData[23359:23328];
//        ram[81856] <= InputData[23391:23360];
//        ram[81857] <= InputData[23423:23392];
//        ram[81858] <= InputData[23455:23424];
//        ram[81859] <= InputData[23487:23456];
//        ram[81860] <= InputData[23519:23488];
//        ram[81861] <= InputData[23551:23520];
//        ram[81862] <= InputData[23583:23552];
//        ram[81863] <= InputData[23615:23584];
//        ram[81864] <= InputData[23647:23616];
//        ram[81865] <= InputData[23679:23648];
//        ram[81866] <= InputData[23711:23680];
//        ram[81867] <= InputData[23743:23712];
//        ram[81868] <= InputData[23775:23744];
//        ram[81869] <= InputData[23807:23776];
//        ram[81870] <= InputData[23839:23808];
//        ram[81871] <= InputData[23871:23840];
//        ram[81872] <= InputData[23903:23872];
//        ram[81873] <= InputData[23935:23904];
//        ram[81874] <= InputData[23967:23936];
//        ram[81875] <= InputData[23999:23968];
//        ram[81876] <= InputData[24031:24000];
//        ram[81877] <= InputData[24063:24032];
//        ram[81878] <= InputData[24095:24064];
//        ram[81879] <= InputData[24127:24096];
//        ram[81880] <= InputData[24159:24128];
//        ram[81881] <= InputData[24191:24160];
//        ram[81882] <= InputData[24223:24192];
//        ram[81883] <= InputData[24255:24224];
//        ram[81884] <= InputData[24287:24256];
//        ram[81885] <= InputData[24319:24288];
//        ram[81886] <= InputData[24351:24320];
//        ram[81887] <= InputData[24383:24352];
//        ram[81888] <= InputData[24415:24384];
//        ram[81889] <= InputData[24447:24416];
//        ram[81890] <= InputData[24479:24448];
//        ram[81891] <= InputData[24511:24480];
//        ram[81892] <= InputData[24543:24512];
//        ram[81893] <= InputData[24575:24544];
//        ram[81894] <= InputData[24607:24576];
//        ram[81895] <= InputData[24639:24608];
//        ram[81896] <= InputData[24671:24640];
//        ram[81897] <= InputData[24703:24672];
//        ram[81898] <= InputData[24735:24704];
//        ram[81899] <= InputData[24767:24736];
//        ram[81900] <= InputData[24799:24768];
//        ram[81901] <= InputData[24831:24800];
//        ram[81902] <= InputData[24863:24832];
//        ram[81903] <= InputData[24895:24864];
//        ram[81904] <= InputData[24927:24896];
//        ram[81905] <= InputData[24959:24928];
//        ram[81906] <= InputData[24991:24960];
//        ram[81907] <= InputData[25023:24992];
//        ram[81908] <= InputData[25055:25024];
//        ram[81909] <= InputData[25087:25056];
//    end

    always @(posedge clk) begin
//        if (rst) begin
//            InputAddr <= 17'd82150;
//            tmp <= InputData;
//        end 
//        else
        begin
            if (InputAddr >= 82150 && InputAddr <= 82933) begin
                ram[InputAddr] <= tmp[DATA_WIDTH-1:0];
                tmp <= {{(32){1'b0}},tmp[25087:32]};
                InputAddr <= InputAddr + 1;
            end
        end
    end
    
//    assign data = ram[addr];
    always @(posedge clk) begin
       if (str)
          ram[addr] <=  MDin;
    end
    
    
    always @(posedge clk or addr) begin
        data <= ram[addr];  //��
    end
          
    
endmodule



`timescale 1ns / 1ps

module test_uart_top();

  reg clk;
  reg rst;
  reg rx;
  wire tx;
  wire parity;
  wire [7:0] SEG,AN;

  test_UART uart_top
  (
    .i_clk_sys(clk), //ϵͳʱ��
    .i_rst_n(rst), //ȫ���첽��λ
    .i_uart_rx(rx), //��������,UART���� 
    .o_uart_tx(tx), //��������,UART���
    .o_ld_parity(parity), //У��λ����LED
    .SEG(SEG),
    .AN(AN)
  ); 

  // ʱ������
  always begin
    #1 clk = ~clk;
  end

  // �����ź�
    initial begin
      clk = 0;
      rst = 0;
      // �ȴ�һ��ʱ�䣬Ȼ���ͷ������ź�
      #100000 rst = 1; //t=10T
      // �ȴ�һ��ʱ���ʼ��������
      #100000 rx = 1; //t=11T
  
      // ģ���������
      $display("Receiving data...");
      // ��ʼ�������� 
      //10101011
      #100000 rx = 0; //210us
      #100000 rx = 1;
      #100000 rx = 1;
      #100000 rx = 0;
      #100000 rx = 1;
      #100000 rx = 0;
      #100000 rx = 1;
      #100000 rx = 0;
      #100000 rx = 1;
      #100000 rx = 1;
      
      #100000 rx = 1;
      
      //01000001
      #100000 rx = 0;
      #100000 rx = 1;
      #100000 rx = 0;
      #100000 rx = 0;
      #100000 rx = 0;
      #100000 rx = 0;
      #100000 rx = 0;
      #100000 rx = 1;
      #100000 rx = 0;
      #100000 rx = 1;
      
      #100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 1;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 0;
#100000 rx = 1;

#100000 rx = 1;

    #6000000; // ���ܺͷ���֮����һ��ʱ�� t=512T
    //��ʼ�������� 
    
    //��������=01000001(0x41)
    #100000  // ��ʼλ t=513T 0
    #100000  // ��һ������λ t=523T 1
    #100000; // �ڶ�������λ t=533T 0
    #100000; // ����������λ t=543T 0
    #100000; // ���ĸ�����λ t=553T 0
    #100000; // ���������λ t=563T 0
    #100000; // ����������λ t=573T 0
    #100000; // ���߸�����λ t=583T 1
    #100000; // �ڰ˸�����λ t=593T 0
    #100000; //ֹͣλ t=603T 1
    
    //��������=01000010(0x42)
    #100000  // ��ʼλ t=613T 0
    #100000  // ��һ������λ t=623T 0
    #100000; // �ڶ�������λ t=633T 1
    #100000; // ����������λ t=643T 0
    #100000; // ���ĸ�����λ t=653T 0
    #100000; // ���������λ t=663T 0
    #100000; // ����������λ t=673T 0
    #100000; // ���߸�����λ t=683T 1
    #100000; // �ڰ˸�����λ t=693T 0
    #100000; //ֹͣλ t=703T 1
    
    //��������=01000011(0x43)
    #100000  // ��ʼλ t=713T 0
    #100000  // ��һ������λ t=723T 1
    #100000; // �ڶ�������λ t=733T 1
    #100000; // ����������λ t=743T 0
    #100000; // ���ĸ�����λ t=753T 0
    #100000; // ���������λ t=763T 0
    #100000; // ����������λ t=773T 0
    #100000; // ���߸�����λ t=783T 1
    #100000; // �ڰ˸�����λ t=793T 0
    #100000; //ֹͣλ t=803T 1
    
    //��������=01000100(0x44)
    #100000  // ��ʼλ t=813T 0
    #100000  // ��һ������λ t=823T 0
    #100000; // �ڶ�������λ t=833T 0
    #100000; // ����������λ t=843T 1
    #100000; // ���ĸ�����λ t=853T 0
    #100000; // ���������λ t=863T 0
    #100000; // ����������λ t=873T 0
    #100000; // ���߸�����λ t=883T 1
    #100000; // �ڰ˸�����λ t=893T 0
    #100000; //ֹͣλ t=903T 1
    
    #1000000; //���ͽ������������һ��ʱ�� t=1003T
      
      $finish; // ��������
    end

endmodule
